library verilog;
use verilog.vl_types.all;
entity CODDOSACUATRO_vlg_vec_tst is
end CODDOSACUATRO_vlg_vec_tst;
