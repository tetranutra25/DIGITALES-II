library verilog;
use verilog.vl_types.all;
entity RelojHoras_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end RelojHoras_vlg_sample_tst;
