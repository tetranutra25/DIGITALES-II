library verilog;
use verilog.vl_types.all;
entity ImplementacionRelojDigital_vlg_sample_tst is
    port(
        CLk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ImplementacionRelojDigital_vlg_sample_tst;
