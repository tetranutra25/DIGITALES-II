library verilog;
use verilog.vl_types.all;
entity ModOchoTruncadoSeis_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ModOchoTruncadoSeis_vlg_sample_tst;
