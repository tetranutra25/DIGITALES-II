library verilog;
use verilog.vl_types.all;
entity CODDOSACUATRO_vlg_check_tst is
    port(
        X               : in     vl_logic;
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CODDOSACUATRO_vlg_check_tst;
