library verilog;
use verilog.vl_types.all;
entity ALUCOMPLETA_vlg_vec_tst is
end ALUCOMPLETA_vlg_vec_tst;
