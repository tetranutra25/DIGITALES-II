library verilog;
use verilog.vl_types.all;
entity CODEDIECISEISACUATRO is
    port(
        A               : out    vl_logic;
        D8              : in     vl_logic;
        D10             : in     vl_logic;
        D9              : in     vl_logic;
        D11             : in     vl_logic;
        D13             : in     vl_logic;
        D12             : in     vl_logic;
        D14             : in     vl_logic;
        D15             : in     vl_logic;
        B               : out    vl_logic;
        D4              : in     vl_logic;
        D6              : in     vl_logic;
        D5              : in     vl_logic;
        D7              : in     vl_logic;
        C               : out    vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        D               : out    vl_logic;
        D1              : in     vl_logic;
        D0              : in     vl_logic
    );
end CODEDIECISEISACUATRO;
