library verilog;
use verilog.vl_types.all;
entity RelojHoras_vlg_vec_tst is
end RelojHoras_vlg_vec_tst;
