library verilog;
use verilog.vl_types.all;
entity FlipFlop_vlg_vec_tst is
end FlipFlop_vlg_vec_tst;
