library verilog;
use verilog.vl_types.all;
entity ModOchoTruncadoCinco_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ModOchoTruncadoCinco_vlg_sample_tst;
