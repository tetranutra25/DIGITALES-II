library verilog;
use verilog.vl_types.all;
entity CODDOSACUATRO is
    port(
        X               : out    vl_logic;
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        Y               : out    vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic
    );
end CODDOSACUATRO;
