library verilog;
use verilog.vl_types.all;
entity COMPRIMIDO_vlg_vec_tst is
end COMPRIMIDO_vlg_vec_tst;
