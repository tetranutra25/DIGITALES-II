library verilog;
use verilog.vl_types.all;
entity CODEDIECISEISACUATRO_vlg_vec_tst is
end CODEDIECISEISACUATRO_vlg_vec_tst;
