library verilog;
use verilog.vl_types.all;
entity ModOcho_vlg_vec_tst is
end ModOcho_vlg_vec_tst;
