library verilog;
use verilog.vl_types.all;
entity BCDaSIETE_vlg_vec_tst is
end BCDaSIETE_vlg_vec_tst;
