library verilog;
use verilog.vl_types.all;
entity COMPRIMIDO_vlg_check_tst is
    port(
        E3              : in     vl_logic;
        E4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end COMPRIMIDO_vlg_check_tst;
