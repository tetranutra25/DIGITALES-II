library verilog;
use verilog.vl_types.all;
entity RelojSegundero_vlg_vec_tst is
end RelojSegundero_vlg_vec_tst;
