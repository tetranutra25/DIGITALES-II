library verilog;
use verilog.vl_types.all;
entity DECOCUATROADIECISEIS_vlg_vec_tst is
end DECOCUATROADIECISEIS_vlg_vec_tst;
