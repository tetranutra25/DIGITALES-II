library verilog;
use verilog.vl_types.all;
entity ModDieciseis_vlg_vec_tst is
end ModDieciseis_vlg_vec_tst;
