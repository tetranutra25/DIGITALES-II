library verilog;
use verilog.vl_types.all;
entity Pruebas_vlg_check_tst is
    port(
        A0              : in     vl_logic;
        B0              : in     vl_logic;
        C0              : in     vl_logic;
        D0              : in     vl_logic;
        E0              : in     vl_logic;
        F0              : in     vl_logic;
        G0              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Pruebas_vlg_check_tst;
