library verilog;
use verilog.vl_types.all;
entity Pruebas is
    port(
        A0              : out    vl_logic;
        C               : in     vl_logic;
        B               : in     vl_logic;
        D               : in     vl_logic;
        A               : in     vl_logic;
        B0              : out    vl_logic;
        C0              : out    vl_logic;
        D0              : out    vl_logic;
        E0              : out    vl_logic;
        F0              : out    vl_logic;
        G0              : out    vl_logic
    );
end Pruebas;
