-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Tue Mar 15 12:21:16 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Pruebas IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		D :  IN  STD_LOGIC;
		A0 :  OUT  STD_LOGIC;
		B0 :  OUT  STD_LOGIC;
		C0 :  OUT  STD_LOGIC;
		D0 :  OUT  STD_LOGIC;
		E0 :  OUT  STD_LOGIC;
		F0 :  OUT  STD_LOGIC;
		G0 :  OUT  STD_LOGIC
	);
END Pruebas;

ARCHITECTURE bdf_type OF Pruebas IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;


BEGIN 



A0 <= C OR SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1 OR A;


SYNTHESIZED_WIRE_0 <= B AND D;


SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59 AND SYNTHESIZED_WIRE_60 AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_38 <= C AND D;


SYNTHESIZED_WIRE_19 <= C AND D;


SYNTHESIZED_WIRE_42 <= C AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_40 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59 AND C;


SYNTHESIZED_WIRE_41 <= A AND SYNTHESIZED_WIRE_60 AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_44 <= B AND SYNTHESIZED_WIRE_60 AND D;


SYNTHESIZED_WIRE_43 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59 AND SYNTHESIZED_WIRE_60 AND SYNTHESIZED_WIRE_61;


B0 <= A OR SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20;


SYNTHESIZED_WIRE_47 <= C AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_45 <= A AND SYNTHESIZED_WIRE_60 AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_46 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59 AND SYNTHESIZED_WIRE_60 AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_50 <= SYNTHESIZED_WIRE_60 AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_48 <= SYNTHESIZED_WIRE_58 AND B AND SYNTHESIZED_WIRE_60;


SYNTHESIZED_WIRE_49 <= B AND C AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_53 <= C AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_58 AND B AND SYNTHESIZED_WIRE_60;


SYNTHESIZED_WIRE_52 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59 AND C;


SYNTHESIZED_WIRE_58 <= NOT(A);



C0 <= B OR SYNTHESIZED_WIRE_38 OR SYNTHESIZED_WIRE_60;


SYNTHESIZED_WIRE_59 <= NOT(B);



SYNTHESIZED_WIRE_60 <= NOT(C);



SYNTHESIZED_WIRE_61 <= NOT(D);



SYNTHESIZED_WIRE_55 <= SYNTHESIZED_WIRE_40 OR SYNTHESIZED_WIRE_41 OR SYNTHESIZED_WIRE_42;


SYNTHESIZED_WIRE_54 <= SYNTHESIZED_WIRE_43 OR SYNTHESIZED_WIRE_44;


E0 <= SYNTHESIZED_WIRE_45 OR SYNTHESIZED_WIRE_46 OR SYNTHESIZED_WIRE_47;


F0 <= A OR SYNTHESIZED_WIRE_48 OR SYNTHESIZED_WIRE_49 OR SYNTHESIZED_WIRE_50;


G0 <= A OR SYNTHESIZED_WIRE_51 OR SYNTHESIZED_WIRE_52 OR SYNTHESIZED_WIRE_53;


D0 <= SYNTHESIZED_WIRE_54 OR SYNTHESIZED_WIRE_55;


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_60 AND SYNTHESIZED_WIRE_61;


END bdf_type;