library verilog;
use verilog.vl_types.all;
entity ModOchoTruncadoSeis_vlg_vec_tst is
end ModOchoTruncadoSeis_vlg_vec_tst;
