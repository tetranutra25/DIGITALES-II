library verilog;
use verilog.vl_types.all;
entity ModDieciseisTruncadoDiez_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ModDieciseisTruncadoDiez_vlg_sample_tst;
