library verilog;
use verilog.vl_types.all;
entity ModDieciseisTruncadoDiez_vlg_vec_tst is
end ModDieciseisTruncadoDiez_vlg_vec_tst;
