library verilog;
use verilog.vl_types.all;
entity ModOchoTruncadoCinco_vlg_vec_tst is
end ModOchoTruncadoCinco_vlg_vec_tst;
