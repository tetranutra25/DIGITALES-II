library verilog;
use verilog.vl_types.all;
entity Pruebas_vlg_vec_tst is
end Pruebas_vlg_vec_tst;
