library verilog;
use verilog.vl_types.all;
entity ImplementacionRelojDigital_vlg_vec_tst is
end ImplementacionRelojDigital_vlg_vec_tst;
