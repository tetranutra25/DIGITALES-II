library verilog;
use verilog.vl_types.all;
entity ModCuatroTruncadoTres_vlg_vec_tst is
end ModCuatroTruncadoTres_vlg_vec_tst;
