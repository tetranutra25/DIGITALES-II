library verilog;
use verilog.vl_types.all;
entity ALUCOMPLETA_vlg_check_tst is
    port(
        C4              : in     vl_logic;
        K0              : in     vl_logic;
        K1              : in     vl_logic;
        K2              : in     vl_logic;
        K3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ALUCOMPLETA_vlg_check_tst;
