library verilog;
use verilog.vl_types.all;
entity ImplementacionRelojDigital_vlg_check_tst is
    port(
        CLK1Hz          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ImplementacionRelojDigital_vlg_check_tst;
